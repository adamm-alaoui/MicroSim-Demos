module simple_logic (
    input a,
    input b,
    input c,
    output out
);

    // Perform a logical OR operation
    assign out = a | b | c;

endmodule
